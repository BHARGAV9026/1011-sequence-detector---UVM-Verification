package pkg;
`include "uvm_macros.svh"
    import uvm_pkg::*;
   
  
  `include "xtn.sv"
  `include "agt_config.sv"
  `include "sequence.sv"
  `include "sequencer.sv"
  `include "driver.sv"
  `include "monitor.sv"
 
  `include "agent.sv"
  `include "sb.sv"
  
  `include "env.sv"
  `include "test.sv"
   
endpackage